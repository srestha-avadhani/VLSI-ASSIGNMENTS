* SPICE3 file created from inverter.ext - technology: scmos

.option scale=0.09u

M1000 Out in gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1001 Out in vdd w_n20_n11# pfet w=25 l=2
+  ad=125 pd=60 as=125 ps=60
C0 w_n20_n11# vdd 0.12fF
C1 w_n20_n11# in 0.08fF
C2 gnd Out 0.10fF
C3 w_n20_n11# Out 0.06fF
C4 in gnd 0.05fF
C5 vdd Out 0.29fF
C6 in Out 0.05fF
C7 gnd Gnd 0.16fF
C8 Out Gnd 0.09fF
C9 vdd Gnd 0.04fF
C10 in Gnd 0.17fF
C11 w_n20_n11# Gnd 1.37fF
