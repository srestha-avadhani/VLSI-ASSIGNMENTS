* SPICE3 file created from ringosc.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale = 0.09u
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

M1 b11 b10 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M2 b11 b10 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M3 b10 b9 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M4 b10 b9 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M5 b12 b11 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M6 b12 b11 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M7 b13 b12 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M8 b13 b12 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M9 b14 b13 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M10 b14 b13 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M11 b15 b14 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M12 b15 b14 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M13 b17 b16 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M14 b17 b16 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M15 b16 b15 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M16 b16 b15 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M17 b18 b17 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M18 b18 b17 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M19 b19 b18 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M20 b19 b18 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M21 b20 b19 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M22 b20 b19 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M23 b21 b20 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M24 b21 b20 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M25 b22 b21 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M26 b22 b21 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M27 b23 b22 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M28 b23 b22 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M29 b24 b23 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M30 b24 b23 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M31 b26 b25 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M32 b26 b25 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M33 b25 b24 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M34 b25 b24 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M35 b27 b26 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M36 b27 b26 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M37 b28 b27 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M38 b28 b27 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M39 b29 b28 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M40 b29 b28 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M41 b30 b29 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M42 b30 b29 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M43 a1 b30 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M44 a1 b30 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M45 b1 a1 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M46 b1 a1 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M47 b2 b1 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M48 b2 b1 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M49 b3 b2 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M50 b3 b2 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M51 b4 b3 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M52 b4 b3 gnd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M53 b5 b4 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M54 b5 b4 gnd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M55 b6 b5 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M56 b6 b5 gnd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M57 b8 b7 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M58 b8 b7 gnd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M59 b7 b6 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M60 b7 b6 gnd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M61 b9 b8 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M62 b9 b8 gnd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60

C0 b10 gnd 0.26fF
C1 vdd b6 0.08fF
C2 b29 b30 0.05fF
C3 b10 gnd 0.26fF
C4 vdd b3 0.29fF
C5 b9 vdd 0.08fF
C6 gnd b20 0.21fF
C7 b5 gnd 0.05fF
C8 gnd b27 0.10fF
C9 b11 b12 0.05fF
C10 vdd vdd 0.12fF
C11 vdd b14 0.06fF
C12 vdd gnd 0.12fF
C13 b25 gnd 0.10fF
C14 gnd b29 0.10fF
C15 gnd a1 0.49fF
C16 vdd b17 0.29fF
C17 vdd gnd 0.12fF
C18 vdd b8 0.06fF
C19 vdd b30 0.29fF
C20 b29 gnd 0.05fF
C21 b30 a1 0.05fF
C22 b10 gnd 0.26fF
C23 vdd vdd 0.12fF
C24 b11 gnd 0.10fF
C25 b7 vdd 0.06fF
C26 gnd b23 0.10fF
C27 b30 vdd 0.08fF
C28 gnd b22 0.10fF
C29 gnd b21 0.10fF
C30 vdd b27 0.08fF
C31 b20 vdd 0.05fF
C32 gnd b14 0.10fF
C33 vdd b10 0.08fF
C34 vdd b26 0.08fF
C35 gnd b19 0.10fF
C36 a1 b1 0.05fF
C37 gnd b28 0.10fF
C38 vdd b24 0.08fF
C39 vdd b26 0.06fF
C40 gnd b4 0.10fF
C41 vdd b29 0.08fF
C42 gnd b18 0.10fF
C43 vdd a1 0.08fF
C44 b7 b8 0.05fF
C45 vdd b25 0.08fF
C46 vdd b24 0.06fF
C47 b28 gnd 0.05fF
C48 vdd b23 0.08fF
C49 b9 vdd 0.06fF
C50 vdd b10 0.06fF
C51 b10 gnd 0.26fF
C52 vdd b6 0.06fF
C53 vdd b22 0.08fF
C54 b10 gnd 0.26fF
C55 vdd b21 0.08fF
C56 vdd b2 0.29fF
C57 gnd b12 0.10fF
C58 vdd vdd 0.12fF
C59 vdd b12 0.29fF
C60 vdd vdd 0.12fF
C61 vdd b19 0.08fF
C62 vdd b1 0.29fF
C63 vdd vdd 0.12fF
C64 b25 b26 0.05fF
C65 b9 gnd 0.05fF
C66 vdd b4 0.08fF
C67 vdd b18 0.08fF
C68 vdd vdd 0.12fF
C69 vdd vdd 0.12fF
C70 gnd b30 0.26fF
C71 vdd vdd 0.12fF
C72 b23 b24 0.05fF
C73 b3 gnd 0.05fF
C74 vdd b17 0.08fF
C75 vdd b29 0.06fF
C76 vdd b13 0.29fF
C77 gnd b30 0.26fF
C78 vdd vdd 0.12fF
C79 b7 b6 0.05fF
C80 b9 b8 0.05fF
C81 b30 vdd 0.04fF
C82 vdd b5 0.06fF
C83 gnd b30 0.26fF
C84 vdd b7 0.08fF
C85 vdd vdd 0.12fF
C86 vdd b12 0.06fF
C87 gnd b30 0.26fF
C88 vdd vdd 0.12fF
C89 b11 b10 0.05fF
C90 b16 gnd 0.10fF
C91 vdd vdd 0.12fF
C92 b20 gnd 0.05fF
C93 b1 gnd 0.05fF
C94 gnd b20 0.21fF
C95 vdd vdd 0.12fF
C96 vdd vdd 0.12fF
C97 vdd b26 0.29fF
C98 gnd b20 0.21fF
C99 vdd gnd 0.12fF
C100 vdd vdd 0.12fF
C101 gnd b20 0.21fF
C102 gnd b17 0.10fF
C103 gnd b8 0.29fF
C104 vdd b24 0.29fF
C105 vdd vdd 0.12fF
C106 b28 b29 0.05fF
C107 b7 gnd 0.29fF
C108 gnd b3 0.10fF
C109 vdd b28 0.08fF
C110 b10 gnd 0.26fF
C111 b5 b6 0.05fF
C112 vdd b3 0.06fF
C113 b12 b13 0.05fF
C114 gnd b2 0.10fF
C115 b10 gnd 0.26fF
C116 b15 gnd 0.05fF
C117 vdd b5 0.08fF
C118 b8 gnd 0.05fF
C119 b11 vdd 0.06fF
C120 vdd b20 0.06fF
C121 gnd b1 0.10fF
C122 gnd b10 0.43fF
C123 gnd b20 0.21fF
C124 vdd b29 0.29fF
C125 vdd a1 0.06fF
C126 b9 gnd 0.29fF
C127 vdd vdd 0.12fF
C128 vdd vdd 0.12fF
C129 vdd vdd 0.12fF
C130 vdd gnd 0.12fF
C131 gnd b6 0.29fF
C132 b2 gnd 0.05fF
C133 b10 gnd 0.26fF
C134 b14 vdd 0.29fF
C135 vdd b2 0.08fF
C136 gnd b16 0.05fF
C137 b15 vdd 0.06fF
C138 b27 gnd 0.05fF
C139 b16 b17 0.05fF
C140 vdd gnd 0.12fF
C141 b20 b21 0.05fF
C142 gnd b15 0.10fF
C143 b10 gnd 0.26fF
C144 b26 gnd 0.05fF
C145 b19 b20 0.05fF
C146 gnd b20 0.21fF
C147 b24 gnd 0.05fF
C148 gnd b26 0.10fF
C149 b6 gnd 0.05fF
C150 b25 gnd 0.05fF
C151 gnd b24 0.10fF
C152 vdd vdd 0.12fF
C153 vdd b4 0.06fF
C154 b13 vdd 0.06fF
C155 b14 vdd 0.08fF
C156 b23 gnd 0.05fF
C157 gnd b14 0.05fF
C158 b4 b5 0.05fF
C159 b22 gnd 0.05fF
C160 vdd b10 0.29fF
C161 b21 gnd 0.05fF
C162 vdd vdd 0.12fF
C163 vdd b16 0.06fF
C164 b12 vdd 0.08fF
C165 vdd vdd 0.12fF
C166 vdd b27 0.06fF
C167 vdd b20 0.29fF
C168 b19 gnd 0.05fF
C169 gnd b20 0.21fF
C170 b18 gnd 0.05fF
C171 gnd b8 0.10fF
C172 b25 vdd 0.06fF
C173 b3 b4 0.05fF
C174 b17 gnd 0.05fF
C175 b13 b14 0.05fF
C176 vdd a1 0.29fF
C177 b7 gnd 0.10fF
C178 vdd b3 0.08fF
C179 vdd vdd 0.12fF
C180 b30 gnd 0.05fF
C181 gnd b5 0.29fF
C182 vdd b23 0.06fF
C183 b15 vdd 0.29fF
C184 vdd b22 0.06fF
C185 vdd b15 0.08fF
C186 vdd b21 0.06fF
C187 b13 vdd 0.08fF
C188 b26 b27 0.05fF
C189 vdd b1 0.08fF
C190 vdd b19 0.06fF
C191 a1 gnd 0.05fF
C192 b13 gnd 0.10fF
C193 vdd b28 0.06fF
C194 gnd b30 0.26fF
C195 b25 b24 0.05fF
C196 gnd b4 0.29fF
C197 vdd b18 0.06fF
C198 gnd b30 0.26fF
C199 b16 b15 0.05fF
C200 b9 gnd 0.10fF
C201 vdd gnd 0.12fF
C202 gnd b30 0.26fF
C203 vdd vdd 0.12fF
C204 vdd vdd 0.12fF
C205 gnd b10 0.05fF
C206 gnd b30 0.26fF
C207 gnd b6 0.10fF
C208 b22 b23 0.05fF
C209 vdd b17 0.06fF
C210 b30 gnd 0.43fF
C211 b12 gnd 0.05fF
C212 gnd b30 0.26fF
C213 b11 gnd 0.05fF
C214 b11 vdd 0.29fF
C215 b21 b22 0.05fF
C216 b9 b10 0.05fF
C217 vdd b2 0.06fF
C218 b13 gnd 0.05fF
C219 vdd b27 0.29fF
C220 b20 gnd 0.35fF
C221 b16 vdd 0.29fF
C222 vdd b8 0.08fF
C223 b4 gnd 0.05fF
C224 gnd b20 0.21fF
C225 b18 b19 0.05fF
C226 vdd b1 0.06fF
C227 b27 b28 0.05fF
C228 b25 vdd 0.29fF
C229 b17 b18 0.05fF
C230 vdd b30 0.06fF
C231 gnd b5 0.10fF
C232 b11 vdd 0.08fF
C233 b7 gnd 0.05fF
C234 vdd b23 0.29fF
C235 b2 b3 0.05fF
C236 vdd b22 0.29fF
C237 vdd b21 0.29fF
C238 b1 b2 0.05fF
C239 b15 b14 0.05fF
C240 b20 vdd 0.08fF
C241 gnd b20 0.21fF
C242 vdd b16 0.08fF
C243 vdd b19 0.29fF
C244 vdd b28 0.29fF
C245 vdd b18 0.29fF
C246 gnd Gnd 0.16fF
C247 gnd Gnd 0.04fF
C248 b8 Gnd 0.29fF
C249 vdd Gnd 1.37fF
C250 gnd Gnd 0.16fF
C251 gnd Gnd 0.04fF
C252 b6 Gnd 0.30fF
C253 vdd Gnd 1.37fF
C254 gnd Gnd 0.16fF
C255 gnd Gnd 0.04fF
C256 b7 Gnd 0.30fF
C257 vdd Gnd 1.37fF
C258 gnd Gnd 0.16fF
C259 gnd Gnd 0.04fF
C260 b5 Gnd 0.30fF
C261 vdd Gnd 1.37fF
C262 gnd Gnd 0.16fF
C263 gnd Gnd 0.04fF
C264 b4 Gnd 0.30fF
C265 vdd Gnd 1.37fF
C266 gnd Gnd 0.16fF
C267 gnd Gnd 0.04fF
C268 b3 Gnd 0.31fF
C269 vdd Gnd 1.37fF
C270 gnd Gnd 0.16fF
C271 vdd Gnd 0.04fF
C272 b2 Gnd 0.31fF
C273 vdd Gnd 1.37fF
C274 gnd Gnd 0.16fF
C275 vdd Gnd 0.04fF
C276 b1 Gnd 0.32fF
C277 vdd Gnd 1.37fF
C278 gnd Gnd 0.16fF
C279 vdd Gnd 0.04fF
C280 a1 Gnd 1.75fF
C281 vdd Gnd 1.37fF
C282 gnd Gnd 0.16fF
C283 vdd Gnd 0.04fF
C284 vdd Gnd 1.37fF
C285 gnd Gnd 0.16fF
C286 b30 Gnd 0.88fF
C287 vdd Gnd 0.04fF
C288 b29 Gnd 0.30fF
C289 vdd Gnd 1.37fF
C290 gnd Gnd 0.16fF
C291 vdd Gnd 0.04fF
C292 b28 Gnd 0.30fF
C293 vdd Gnd 1.37fF
C294 gnd Gnd 0.16fF
C295 vdd Gnd 0.04fF
C296 b27 Gnd 0.30fF
C297 vdd Gnd 1.37fF
C298 gnd Gnd 0.16fF
C299 vdd Gnd 0.04fF
C300 b26 Gnd 0.29fF
C301 vdd Gnd 1.37fF
*C302 gnd Gnd 0.16fF
C303 vdd Gnd 0.04fF
C304 b24 Gnd 0.29fF
C305 vdd Gnd 1.37fF
*C306 gnd Gnd 0.16fF
C307 vdd Gnd 0.04fF
C308 b25 Gnd 0.29fF
C309 vdd Gnd 1.37fF
*C310 gnd Gnd 0.16fF
C311 vdd Gnd 0.04fF
C312 b23 Gnd 0.29fF
C313 vdd Gnd 1.37fF
*C314 gnd Gnd 0.16fF
C315 vdd Gnd 0.04fF
C316 b22 Gnd 0.30fF
C317 vdd Gnd 1.37fF
*C318 gnd Gnd 0.16fF
C319 vdd Gnd 0.04fF
C320 b21 Gnd 0.30fF
C321 vdd Gnd 1.37fF
*C322 gnd Gnd 0.16fF
C323 vdd Gnd 0.04fF
C324 vdd Gnd 1.37fF
*C325 gnd Gnd 0.16fF
C326 b20 Gnd 0.94fF
C327 vdd Gnd 0.04fF
C328 b19 Gnd 0.29fF
C329 vdd Gnd 1.37fF
*C330 gnd Gnd 0.16fF
C331 vdd Gnd 0.04fF
C332 b18 Gnd 0.30fF
C333 vdd Gnd 1.37fF
*C334 gnd Gnd 0.16fF
C335 vdd Gnd 0.04fF
C336 b17 Gnd 0.29fF
C337 vdd Gnd 1.37fF
*C338 gnd Gnd 0.16fF
C339 vdd Gnd 0.04fF
C340 b15 Gnd 0.30fF
C341 vdd Gnd 1.37fF
*C342 gnd Gnd 0.16fF
C343 vdd Gnd 0.04fF
C344 b16 Gnd 0.30fF
C345 vdd Gnd 1.37fF
*C346 gnd Gnd 0.16fF
C347 vdd Gnd 0.04fF
C348 b14 Gnd 0.29fF
C349 vdd Gnd 1.37fF
*C350 gnd Gnd 0.16fF
C351 vdd Gnd 0.04fF
C352 b13 Gnd 0.29fF
C353 vdd Gnd 1.37fF
C355 vdd Gnd 0.04fF
C356 b12 Gnd 0.29fF
C357 vdd Gnd 1.37fF
*C358 gnd Gnd 0.16fF
C359 vdd Gnd 0.04fF
C360 b11 Gnd 0.30fF
C361 vdd Gnd 1.37fF
*C362 gnd Gnd 0.16fF
C363 b10 Gnd 2.39fF
C364 vdd Gnd 0.04fF
C365 b9 Gnd 0.29fF
C366 vdd Gnd 1.37fF
*C367 gnd Gnd 0.16fF
C368 vdd Gnd 0.04fF
C369 vdd Gnd 1.37fF

.tran 0.1n 200n

.ic v(a1) = 1.8

.measure tran tperiod
+ TRIG v(a1) VAL='SUPPLY/2' RISE=1
+ TARG v(a1) VAL='SUPPLY/2' RISE=2

.measure tran tpdr
+ TRIG v(b1) VAL='SUPPLY/2' FALL=1
+ TARG v(b2) VAL='SUPPLY/2' RISE=1

.measure tran tpdf
+ TRIG v(b1) VAL='SUPPLY/2' RISE=1
+ TARG v(b2) VAL='SUPPLY/2' FALL=1

.measure tran tpd param='(tpdr+tpdf)/2' goal=0

.control

run

.endc
