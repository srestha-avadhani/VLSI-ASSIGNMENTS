magic
tech scmos
timestamp 1613411443
<< nwell >>
rect -20 -11 11 33
<< ntransistor >>
rect -6 -29 -4 -19
<< ptransistor >>
rect -6 -3 -4 22
<< ndiffusion >>
rect -7 -29 -6 -19
rect -4 -29 -3 -19
<< pdiffusion >>
rect -7 -3 -6 22
rect -4 -3 -3 22
<< ndcontact >>
rect -11 -29 -7 -19
rect -3 -29 1 -19
<< pdcontact >>
rect -11 -3 -7 22
rect -3 -3 1 22
<< polysilicon >>
rect -6 22 -4 25
rect -6 -19 -4 -3
rect -6 -34 -4 -29
<< polycontact >>
rect -10 -16 -6 -12
<< metal1 >>
rect -20 28 11 33
rect -11 22 -7 28
rect -3 -12 1 -3
rect -23 -16 -10 -12
rect -3 -16 17 -12
rect -3 -19 1 -16
rect -11 -37 -7 -29
rect -21 -42 10 -37
<< labels >>
rlabel metal1 -20 28 11 33 5 vdd
rlabel metal1 1 -16 17 -12 1 Out
rlabel metal1 -23 -16 -10 -12 1 in
rlabel metal1 -21 -42 10 -37 1 gnd
<< end >>
